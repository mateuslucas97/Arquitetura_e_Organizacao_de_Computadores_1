library verilog;
use verilog.vl_types.all;
entity func1 is
    port(
        I0              : in     vl_logic;
        I1              : in     vl_logic;
        S               : in     vl_logic;
        \out\           : out    vl_logic
    );
end func1;
