library verilog;
use verilog.vl_types.all;
entity multiplicador is
    port(
        a               : in     vl_logic_vector(7 downto 0);
        b               : in     vl_logic_vector(7 downto 0);
        resultado       : out    vl_logic_vector(7 downto 0)
    );
end multiplicador;
